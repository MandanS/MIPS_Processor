`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Mandan Sharma 
// 
// Create Date:    19:40:08 12/05/2017 
// Design Name: 
// Module Name:    Tile_generator 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Tile_generator(
	input wire clk,
   input wire [9:0] pixel_x,
	input wire [9:0] pixel_y, 
	output wire [13:0] addr_b,
	input wire [15:0] din_b,
	output reg [2:0] Red,Green,
	output reg [1:0] Blue,
	input wire video_on
    );

	 

	 assign addr_b = (pixel_y[8:4] << 5 + pixel_x[9:3]) << 1 ;

		

	// signal declaton

	reg [10:0] addr_reg ;
	reg [7:0] data;
	
	always @(posedge clk) 
		addr_reg <= {din_b[6:0],pixel_y[3:0]};
	


	always @*
	case (addr_reg)
		//code x41 blank letter A
		11'h410 : data = 8'b00000000;
		11'h411 : data = 8'b00000000;
		11'h412 : data = 8'b00111000;
		11'h413 : data = 8'b01101100;
		11'h414 : data = 8'b11000110;
		11'h415 : data = 8'b11000110;
		11'h416 : data = 8'b11000110;
		11'h417 : data = 8'b11111110;
		11'h418 : data = 8'b11000110;
		11'h419 : data = 8'b11000110;
		11'h41A : data = 8'b11000110;
		11'h41B : data = 8'b11000110;
		11'h41C : data = 8'b00000000;
		11'h41D : data = 8'b00000000;
		11'h41E : data = 8'b00000000;
		11'h41F : data = 8'b00000000;
		
		//code x42 blank letter B
	endcase	
		
		
		always@(pixel_x)

		if((video_on && data[pixel_x[2:0]] )== 1'b1)	
					{Red,Green,Blue} = din_b[15:8];
		else				
					{Red,Green,Blue} = 8'h00;

		
		
		
		
		
//initial
//		begin
//		
//		rom_A = {
//
//							8'b00000000,
//							8'b00000000,
//							8'b00111000,
//							8'b01101100,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11111110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_B = {   
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b11111100,
//							8'b01100110,
//							8'b01100110,
//							8'b01100110,
//							8'b01111100,
//							8'b01100110,
//							8'b01100110,
//							8'b01100110,
//							8'b01100110,
//							8'b11111100,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_C = {
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b01111100,
//							8'b11000110,
//							8'b11000110,
//							8'b11000000,
//							8'b11000000,
//							8'b11000000,
//							8'b11000000,
//							8'b11000110,
//							8'b11000110,
//							8'b01111100,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_D = {                            
//							8'b00000000,
//							8'b00000000,
//							8'b11111100,
//							8'b01100110,
//							8'b01100110,
//							8'b01100110,
//							8'b01100110,
//							8'b01100110,
//							8'b01100110,
//							8'b01100110,
//							8'b01100110,
//							8'b11111100,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_E = {
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b11111110,
//							8'b01100110,
//							8'b01100010,
//							8'b01101000,
//							8'b01111000,
//							8'b01111000,
//							8'b01101000,
//							8'b01100010,
//							8'b01100110,
//							8'b11111110,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_F = {    
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b11111110,
//							8'b01100110,
//							8'b01100010,
//							8'b01101000,
//							8'b01111000,
//							8'b01111000,
//							8'b01101000,
//							8'b01100000,
//							8'b01100000,
//							8'b11110000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_G = {  
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b01111100,
//							8'b11000110,
//							8'b11000110,
//							8'b11000000,
//							8'b11000000,
//							8'b11001110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b01111110,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_H = {
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11111110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_I = {    
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b00111100,
//							8'b00011000,
//							8'b00011000,
//							8'b00011000,
//							8'b00011000,
//							8'b00011000,
//							8'b00011000,
//							8'b00011000,
//							8'b00011000,
//							8'b00111100,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_J = {    
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b00011110,
//							8'b00001100,
//							8'b00001100,
//							8'b00001100,
//							8'b00001100,
//							8'b00001100,
//							8'b11001100,
//							8'b11001100,
//							8'b11001100,
//							8'b01111000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_K = {  
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b11100110,
//							8'b01100110,
//							8'b01100110,
//							8'b01101100,
//							8'b01111000,
//							8'b01111000,
//							8'b01101100,
//							8'b01100110,
//							8'b01100110,
//							8'b11100110,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_L = {  
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b11110000,
//							8'b01100000,
//							8'b01100000,
//							8'b01100000,
//							8'b01100000,
//							8'b01100000,
//							8'b01100000,
//							8'b01100010,
//							8'b01100110,
//							8'b11111110,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_M = {    
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b10000010,
//							8'b11000110,
//							8'b11101110,
//							8'b11111110,
//							8'b11111110,
//							8'b11010110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_N = {   
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b10000110,
//							8'b11000110,
//							8'b11100110,
//							8'b11110110,
//							8'b11111110,
//							8'b11011110,
//							8'b11001110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_O = {    
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b01111100,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b01111100,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_P = {    
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b11111100,
//							8'b01100110,
//							8'b01100110,
//							8'b01100110,
//							8'b01100110,
//							8'b01111100,
//							8'b01100000,
//							8'b01100000,
//							8'b01100000,
//							8'b11110000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_Q = {  
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b01111100,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11010110,
//							8'b11011110,
//							8'b01111100,
//							8'b00000110,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_R = {  
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b11111100,
//							8'b01100110,
//							8'b01100110,
//							8'b01100110,
//							8'b01100110,
//							8'b01111100,
//							8'b01101100,
//							8'b01100110,
//							8'b01100110,
//							8'b11100110,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_S = {   
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b01111100,
//							8'b11000110,
//							8'b11000110,
//							8'b01100000,
//							8'b00111000,
//							8'b00001100,
//							8'b00000110,
//							8'b11000110,
//							8'b11000110,
//							8'b01111100,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_T = {   
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b01111110,
//							8'b01111110,
//							8'b01011010,
//							8'b00011000,
//							8'b00011000,
//							8'b00011000,
//							8'b00011000,
//							8'b00011000,
//							8'b00011000,
//							8'b00111100,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_U = {   
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b01111100,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_V = {  
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b01101100,
//							8'b00111000,
//							8'b00010000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_W = {   
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11000110,
//							8'b11010110,
//							8'b11111110,
//							8'b11101110,
//							8'b11000110,
//							8'b10000010,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_X = {    
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b11000110,
//							8'b11000110,
//							8'b01101100,
//							8'b01111100,
//							8'b00111000,
//							8'b00111000,
//							8'b01111100,
//							8'b01101100,
//							8'b11000110,
//							8'b11000110,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_Y = {   
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b01100110,
//							8'b01100110,
//							8'b01100110,
//							8'b01100110,
//							8'b00111100,
//							8'b00011000,
//							8'b00011000,
//							8'b00011000,
//							8'b00011000,
//							8'b00111100,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	                        
//	};                      
//	                        
//		rom_Z = {   
//                            
//							8'b00000000,
//							8'b00000000,
//							8'b11111110,
//							8'b11000110,
//							8'b10000110,
//							8'b00001100,
//							8'b00011000,
//							8'b00110000,
//							8'b01100000,
//							8'b11000010,
//							8'b11000110,
//							8'b11111110,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000,
//							8'b00000000
//	
//	};
//	
//				rom_white = {
//
//	8'hFF,
//	8'hFF,
//	8'hFF,
//	8'hFF,
//	8'hFF,
//	8'hFF,
//	8'hFF,
//	8'hFF,
//	8'hFF,
//	8'hFF,
//	8'hFF,
//	8'hFF,
//	8'hFF,
//	8'hFF,
//	8'hFF,
//	8'hFF
//	
//	};
//	
	
//	
//	end
//	
//	reg [7:0]px;
//
//	
//	always @(din_b[7:0] or pixel_y[3:0])
//		begin
//			case (din_b[7:0])
//
//				8'h41:  px  =  rom_A[din_b];  //  A 
//				8'h42:  px  =  rom_B[din_b[15:0]];  //  B 
//				8'h43:  px  =  rom_C[din_b[15:0]];  //  C 
//				8'h44:  px  =  rom_D[din_b[15:0]];  //  D 
//				8'h45:  px  =  rom_E[din_b[15:0]];  //  E 
//				8'h46:  px  =  rom_F[din_b[15:0]];  //  F 
//				8'h46:  px  =  rom_G[din_b[15:0]];  //  G 
//				8'h48:  px  =  rom_H[din_b[15:0]];  //  H 
//				8'h49:  px  =  rom_I[din_b[15:0]];  //  I 
//				8'h4A:  px  =  rom_J[din_b[15:0]];  //  J 
//				8'h4B:  px  =  rom_K[din_b[15:0]];  //  K 
//				8'h4C:  px  =  rom_L[din_b[15:0]];  //  L 
//				8'h4D:  px  =  rom_M[din_b[15:0]];  //  M 
//				8'h4E:  px  =  rom_N[din_b[15:0]];  //  N 
//				8'h4F:  px  =  rom_O[din_b[15:0]];  //  O 
//				8'h50:  px  =  rom_P[din_b[15:0]];  //  P 
//				8'h51:  px  =  rom_Q[din_b[15:0]];  //  Q 
//				8'h52:  px  =  rom_R[din_b[15:0]];  //  R 
//				8'h53:  px  =  rom_S[din_b[15:0]];  //  S 
//				8'h54:  px  =  rom_T[din_b[15:0]];  //  T 
//				8'h55:  px  =  rom_U[din_b[15:0]];  //  U 
//				8'h56:  px  =  rom_V[din_b[15:0]];  //  V 
//				8'h57:  px  =  rom_W[din_b[15:0]];  //  W 
//				8'h58:  px  =  rom_X[din_b[15:0]];  //  X 
//				8'h59:  px  =  rom_Y[din_b[15:0]];  //  Y 
//				8'h5A:  px  =  rom_Z[din_b[15:0]];  //  Z 
//	
//				default:px =  rom_white[din_b[15:0]];
//			endcase
//		end

	

	

endmodule
